//      // verilator_coverage annotation
        //========================================================================
        // Verilog Components: Registers
        //========================================================================
        
        // Note that we place the register output earlier in the port list since
        // this is one place we might actually want to use positional port
        // binding like this:
        //
        //  logic [p_nbits-1:0] result_B;
        //  vc_Reg#(p_nbits) result_AB( clk, result_B, result_A );
        
        `ifndef VC_REGS_V
        `define VC_REGS_V
        
        //------------------------------------------------------------------------
        // Postive-edge triggered flip-flop
        //------------------------------------------------------------------------
        
        module vc_Reg
        #(
          parameter p_nbits = 1
        )(
 134680   input  logic               clk, // Clock input
 000576   output logic [p_nbits-1:0] q,   // Data output
 000576   input  logic [p_nbits-1:0] d    // Data input
        );
        
 067254   always_ff @( posedge clk )
 067254     q <= d;
        
        endmodule
        
        //------------------------------------------------------------------------
        // Postive-edge triggered flip-flop with reset
        //------------------------------------------------------------------------
        
        module vc_ResetReg
        #(
          parameter p_nbits       = 1,
          parameter p_reset_value = 0
        )(
 202020   input  logic               clk,   // Clock input
 000258   input  logic               reset, // Sync reset input
 014854   output logic [p_nbits-1:0] q,     // Data output
 014872   input  logic [p_nbits-1:0] d      // Data input
        );
        
 100881   always_ff @( posedge clk )
 100881     q <= reset ? p_reset_value : d;
        
        endmodule
        
        //------------------------------------------------------------------------
        // Postive-edge triggered flip-flop with enable
        //------------------------------------------------------------------------
        
        module vc_EnReg
        #(
          parameter p_nbits = 1
        )(
 061129   input  logic               clk,   // Clock input
 000043   input  logic               reset, // Sync reset input
 000809   output logic [p_nbits-1:0] q,     // Data output
 002214   input  logic [p_nbits-1:0] d,     // Data input
 000062   input  logic               en     // Enable input
        );
        
 030543   always_ff @( posedge clk )
 000031     if ( en )
 000031       q <= d;
        
          // Assertions
        
          `ifndef SYNTHESIS
        
          /*
          always_ff @( posedge clk )
            if ( !reset )
              `VC_ASSERT_NOT_X( en );
          */
        
          `endif /* SYNTHESIS */
        
        endmodule
        
        //------------------------------------------------------------------------
        // Postive-edge triggered flip-flop with enable and reset
        //------------------------------------------------------------------------
        
        module vc_EnResetReg
        #(
          parameter p_nbits       = 1,
          parameter p_reset_value = 0
        )(
 000250   input  logic               clk,   // Clock input
 000002   input  logic               reset, // Sync reset input
%000000   output logic [p_nbits-1:0] q,     // Data output
%000000   input  logic [p_nbits-1:0] d,     // Data input
 000004   input  logic               en     // Enable input
        );
        
 000124   always_ff @( posedge clk )
 000022     if ( reset || en )
 000102       q <= reset ? p_reset_value : d;
        
          // Assertions
        
          `ifndef SYNTHESIS
        
          /*
          always_ff @( posedge clk )
            if ( !reset )
              `VC_ASSERT_NOT_X( en );
          */
        
          `endif /* SYNTHESIS */
        
        endmodule
        
        `endif /* VC_REGS_V */
        
        
