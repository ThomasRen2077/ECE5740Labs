//      // verilator_coverage annotation
        //========================================================================
        // Verilog Components: Drop Unit
        //========================================================================
        // Drop unit allows dropping a packet when the drop signal is high. This
        // is useful especially in pipelined processor, when a squash should drop
        // a late arriving memory response.
        
        `ifndef LAB2_PROC_DROP_UNIT_V
        `define LAB2_PROC_DROP_UNIT_V
        
        module lab2_proc_DropUnit
        #(
          parameter p_msg_nbits = 1
        )
        (
 029070   input  logic                   clk,
 000080   input  logic                   reset,
        
          // the drop signal will drop the next arriving packet
        
 000532   input  logic                   drop,
        
 001412   input  logic [p_msg_nbits-1:0] istream_msg,
 008661   input  logic                   istream_val,
 009055   output logic                   istream_rdy,
        
 001412   output logic [p_msg_nbits-1:0] ostream_msg,
 008405   output logic                   ostream_val,
 009147   input  logic                   ostream_rdy
        );
        
          localparam c_state_pass = 1'b0;
          localparam c_state_drop = 1'b1;
        
 000248   logic state;
 000248   logic next_state;
 009159   logic istream_go;
        
          assign istream_go = istream_rdy && istream_val;
        
          // assign output message same as input message
        
          assign ostream_msg = istream_msg;
        
          // next state
        
%000000   always_comb begin
 000151     if ( state == c_state_pass ) begin
        
              // we only go to drop state if there is a drop request and we cannot
              // drop it right away (!istream_en)
 000372       if ( drop && !istream_go )
 000372         next_state = c_state_drop;
              else
 042820         next_state = c_state_pass;
        
 000151     end else begin
        
              // if we are in the drop mode and a message arrives, we can go back
              // to pass state
 000081       if ( istream_go )
 000372         next_state = c_state_pass;
              else
 000081         next_state = c_state_drop;
        
            end
          end
        
          // state outputs
        
%000000   always_comb begin
 000151     if ( state == c_state_pass ) begin
        
              // we combinationally take care of dropping if the packet is already
              // available
 014344       ostream_val = istream_val && !drop;
 014344       istream_rdy  = ostream_rdy;
        
 000151     end else begin
        
              // we just drop the packet
 000151       ostream_val = 1'b0;
 000151       istream_rdy  = 1'b1;
        
            end
          end
        
          // state transitions
        
 014495   always_ff @( posedge clk ) begin
        
 001040     if ( reset )
 001040       state <= c_state_pass;
            else
 013455       state <= next_state;
        
          end
        
        endmodule
        
        `endif /* LAB2_PROC_DROP_UNIT_V */
        
        
