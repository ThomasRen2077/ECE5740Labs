//      // verilator_coverage annotation
        //========================================================================
        // Verilog Components: Arithmetic Components
        //========================================================================
        
        `ifndef VC_ARITHMETIC_V
        `define VC_ARITHMETIC_V
        
        //------------------------------------------------------------------------
        // Adders
        //------------------------------------------------------------------------
        
        module vc_Adder
        #(
          parameter p_nbits = 1
        )(
 000041   input  logic [p_nbits-1:0] in0,
 000664   input  logic [p_nbits-1:0] in1,
%000000   input  logic               cin,
 000359   output logic [p_nbits-1:0] out,
 000980   output logic               cout
        );
        
          // We need to convert cin into a 32-bit value to
          // avoid verilator warnings
        
          assign {cout,out} = in0 + in1 + {{(p_nbits-1){1'b0}},cin};
        
        endmodule
        
        module vc_SimpleAdder
        #(
          parameter p_nbits = 1
        )(
 000016   input  logic [p_nbits-1:0] in0,
 000002   input  logic [p_nbits-1:0] in1,
 000016   output logic [p_nbits-1:0] out
        );
        
          assign out = in0 + in1;
        
        endmodule
        
        //------------------------------------------------------------------------
        // Subtractor
        //------------------------------------------------------------------------
        
        module vc_Subtractor
        #(
          parameter p_nbits = 1
        )(
          input  logic [p_nbits-1:0] in0,
          input  logic [p_nbits-1:0] in1,
          output logic [p_nbits-1:0] out
        );
        
          assign out = in0 - in1;
        
        endmodule
        
        //------------------------------------------------------------------------
        // Incrementer
        //------------------------------------------------------------------------
        
        module vc_Incrementer
        #(
          parameter p_nbits     = 1,
          parameter p_inc_value = 1
        )(
 000082   input  logic [p_nbits-1:0] in,
 000010   output logic [p_nbits-1:0] out
        );
        
          assign out = in + p_inc_value;
        
        endmodule
        
        //------------------------------------------------------------------------
        // ZeroExtender
        //------------------------------------------------------------------------
        
        module vc_ZeroExtender
        #(
          parameter p_in_nbits  = 1,
          parameter p_out_nbits = 8
        )(
          input  logic [p_in_nbits-1:0]  in,
          output logic [p_out_nbits-1:0] out
        );
        
          assign out = { {( p_out_nbits - p_in_nbits ){1'b0}}, in };
        
        endmodule
        
        //------------------------------------------------------------------------
        // SignExtender
        //------------------------------------------------------------------------
        
        module vc_SignExtender
        #(
         parameter p_in_nbits = 1,
         parameter p_out_nbits = 8
        )
        (
          input  logic [p_in_nbits-1:0]  in,
          output logic [p_out_nbits-1:0] out
        );
        
          assign out = { {(p_out_nbits-p_in_nbits){in[p_in_nbits-1]}}, in };
        
        endmodule
        
        //------------------------------------------------------------------------
        // ZeroComparator
        //------------------------------------------------------------------------
        
        module vc_ZeroComparator
        #(
          parameter p_nbits = 1
        )(
 000468   input  logic [p_nbits-1:0] in,
 001866   output logic               out
        );
        
          assign out = ( in == {p_nbits{1'b0}} );
        
        endmodule
        
        //------------------------------------------------------------------------
        // EqComparator
        //------------------------------------------------------------------------
        
        module vc_EqComparator
        #(
          parameter p_nbits = 1
        )(
 000016   input  logic [p_nbits-1:0] in0,
 000468   input  logic [p_nbits-1:0] in1,
 003306   output logic               out
        );
        
          assign out = ( in0 == in1 );
        
        endmodule
        
        //------------------------------------------------------------------------
        // LtComparator
        //------------------------------------------------------------------------
        
        module vc_LtComparator
        #(
          parameter p_nbits = 1
        )(
          input  logic [p_nbits-1:0] in0,
          input  logic [p_nbits-1:0] in1,
          output logic               out
        );
        
          assign out = ( in0 < in1 );
        
        endmodule
        
        //------------------------------------------------------------------------
        // GtComparator
        //------------------------------------------------------------------------
        
        module vc_GtComparator
        #(
          parameter p_nbits = 1
        )(
          input  logic [p_nbits-1:0] in0,
          input  logic [p_nbits-1:0] in1,
          output logic               out
        );
        
          assign out = ( in0 > in1 );
        
        endmodule
        
        //------------------------------------------------------------------------
        // LeftLogicalShifter
        //------------------------------------------------------------------------
        
        module vc_LeftLogicalShifter
        #(
          parameter p_nbits       = 1,
          parameter p_shamt_nbits = 1 )
        (
 000016   input  logic       [p_nbits-1:0] in,
 000126   input  logic [p_shamt_nbits-1:0] shamt,
 000210   output logic       [p_nbits-1:0] out
        );
        
          assign out = ( in << shamt );
        
        endmodule
        
        //------------------------------------------------------------------------
        // RightLogicalShifter
        //------------------------------------------------------------------------
        
        module vc_RightLogicalShifter
        #(
          parameter p_nbits       = 1,
          parameter p_shamt_nbits = 1
        )(
 000468   input  logic       [p_nbits-1:0] in,
 000126   input  logic [p_shamt_nbits-1:0] shamt,
 000480   output logic       [p_nbits-1:0] out
        );
        
          assign out = ( in >> shamt );
        
        endmodule
        
        `endif /* VC_ARITHMETIC_V */
        
        
